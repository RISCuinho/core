`define PAUSE_CLOCK_COUNTER_LIMIT 10
